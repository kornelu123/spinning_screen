module top(
  input btn_0,
  output led_0
);

assign led_0 = btn_0;

endmodule
